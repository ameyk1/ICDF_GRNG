module ROM_coef(clk,rst,		// I: Global IO (clock, reset) 
			  en_coef,      // I: Module Enable signal
			  segment,    	// I: [6:0] Segment (Offset + ROM_trans)
			  coef0,        // O: [20:0] Coefficient 0
			  coef1,        // O: [17:0] Coefficient 1
			  coef2			// O: [17:0] Coefficient 2
			  );

input clk,rst;				// I: Global IO (clock, reset) 
input en_coef;      		// I: Module Enable signal
input [6:0]segment;    		// I: [6:0] Segment (Offset + ROM_trans)
output reg signed [20:0] coef0;	// O: [20:0] Coefficient 0
output reg signed [17:0] coef1;	// O: [17:0] Coefficient 1
output reg signed [17:0] coef2;	// O: [17:0] Coefficient 2

reg [56:0] coef_acc;

always@(*)
	case(segment)
		7'd0 : coef_acc =   57'b0011_11111110101100101___1011_11111010101100___001_000001101001110110;
		7'd1 : coef_acc =   57'b0011_11111111010110110___1011_11110001011100___001_000011110100111000;
		7'd2 : coef_acc =   57'b0011_11111111100100111___1011_11101001000011___001_000101111001110111;
		7'd3 : coef_acc =   57'b0011_11111111101011111___1011_11100000111001___001_000111111110000101;
		7'd4 : coef_acc =   57'b0011_11111111110000001___1011_11011000110101___001_001010000010100100;
		7'd5 : coef_acc =   57'b0011_11111111110010111___1011_11010000110011___001_001100000111101101;
		7'd6 : coef_acc =   57'b0011_11111111110100111___1011_11001000110011___001_001110001101100111;
		7'd7 : coef_acc =   57'b0011_11111111110110011___1011_11000000110100___001_010000010100011000;
		7'd8 : coef_acc =   57'b0011_11111111110111101___1011_10111000110110___001_010010011100000011;
		7'd9 : coef_acc =   57'b0011_11111111111000100___1011_10110000111000___001_010100100100101001;
		7'd10 : coef_acc =   57'b0011_11111111111001010___1011_10101000111010___001_010110101110001100;
		7'd11 : coef_acc =   57'b0011_11111111111001111___1011_10100000111101___001_011000111000101011;
		7'd12 : coef_acc =   57'b0011_11111111111010100___1011_10011001000000___001_011011000100001000;
		7'd13 : coef_acc =   57'b0011_11111111111010111___1011_10010001000011___001_011101010000100011;
		7'd14 : coef_acc =   57'b0011_11111111111011010___1011_10001001000110___001_011111011101111011;
		7'd15 : coef_acc =   57'b0011_11111111111011101___1011_10000001001001___001_100001101100010010;
		7'd16 : coef_acc =   57'b0011_11111111111100000___1011_01111001001101___001_100011111011100111;
		7'd17 : coef_acc =   57'b0011_11111111111100010___1011_01110001010000___001_100110001011111011;
		7'd18 : coef_acc =   57'b0011_11111111111100100___1011_01101001010100___001_101000011101001101;
		7'd19 : coef_acc =   57'b0011_11111111111100101___1011_01100001010111___001_101010101111011110;
		7'd20 : coef_acc =   57'b0011_11111111111100111___1011_01011001011011___001_101101000010101101;
		7'd21 : coef_acc =   57'b0011_11111111111101000___1011_01010001011110___001_101111010110111100;
		7'd22 : coef_acc =   57'b0011_11111111111101010___1011_01001001100010___001_110001101100001000;
		7'd23 : coef_acc =   57'b0011_11111111111101011___1011_01000001100110___001_110100000010010100;
		7'd24 : coef_acc =   57'b0011_11111111111101100___1011_00111001101001___001_110110011001011111;
		7'd25 : coef_acc =   57'b0011_11111111111101101___1011_00110001101101___001_111000110001101000;
		7'd26 : coef_acc =   57'b0011_11111111111101110___1011_00101001110001___001_111011001010110000;
		7'd27 : coef_acc =   57'b0011_11111111111101111___1011_00100001110100___001_111101100100111000;
		7'd28 : coef_acc =   57'b0011_11111111111101111___1011_00011001111000___001_111111111111111110;
		7'd29 : coef_acc =   57'b0011_11111111111110000___1011_00010001111100___010_000010011100000010;
		7'd30 : coef_acc =   57'b0011_11111111111110001___1011_00001010000000___010_000100111001000110;
		7'd31 : coef_acc =   57'b0011_11111111111110001___1011_00000010000100___010_000111010111001001;
		7'd32 : coef_acc =   57'b0011_11111111111110010___1010_11111010000111___010_001001110110001011;
		7'd33 : coef_acc =   57'b0011_11111111111110011___1010_11110010001011___010_001100010110001011;
		7'd34 : coef_acc =   57'b0011_11111111111110011___1010_11101010001111___010_001110110111001011;
		7'd35 : coef_acc =   57'b0011_11111111111110100___1010_11100010010011___010_010001011001001001;
		7'd36 : coef_acc =   57'b0011_11111111111110100___1010_11011010010111___010_010011111100000111;
		7'd37 : coef_acc =   57'b0011_11111111111110101___1010_11010010011011___010_010110100000000011;
		7'd38 : coef_acc =   57'b0011_11111111111110101___1010_11001010011110___010_011001000100111111;
		7'd39 : coef_acc =   57'b0011_11111111111110101___1010_11000010100010___010_011011101010111001;
		7'd40 : coef_acc =   57'b0011_11111111111110110___1010_10111010100110___010_011110010001110010;
		7'd41 : coef_acc =   57'b0011_11111111111110110___1010_10110010101010___010_100000111001101010;
		7'd42 : coef_acc =   57'b0011_11111111111110110___1010_10101010101110___010_100011100010100010;
		7'd43 : coef_acc =   57'b0011_11111111111110111___1010_10100010110010___010_100110001100011000;
		7'd44 : coef_acc =   57'b0011_11111111111110111___1010_10011010110110___010_101000110111001101;
		7'd45 : coef_acc =   57'b0011_11111111111110111___1010_10010010111010___010_101011100011000001;
		7'd46 : coef_acc =   57'b0011_11111111111111000___1010_10001010111101___010_101110001111110101;
		7'd47 : coef_acc =   57'b0011_11111111111111000___1010_10000011000001___010_110000111101100111;
		7'd48 : coef_acc =   57'b0011_11111111111111000___1010_01111011000101___010_110011101100011000;
		7'd49 : coef_acc =   57'b0011_11111111111111000___1010_01110011001001___010_110110011100001000;
		7'd50 : coef_acc =   57'b0011_11111111111111000___1010_01101011001101___010_111001001100110111;
		7'd51 : coef_acc =   57'b0011_11111111111111001___1010_01100011010001___010_111011111110100101;
		7'd52 : coef_acc =   57'b0011_11111111111111001___1010_01011011010101___010_111110110001010010;
		7'd53 : coef_acc =   57'b0011_11111111111111001___1010_01010011011001___0011_000001100100111110;
		7'd54 : coef_acc =   57'b0011_11111111111111001___1010_01001011011101___0011_000100011001101001;
		7'd55 : coef_acc =   57'b0011_11111111111111001___1010_01000011100001___0011_000111001111010100;
		7'd56 : coef_acc =   57'b0011_11111111111111010___1010_00111011100101___0011_001010000101111101;
		7'd57 : coef_acc =   57'b0011_11111111111111010___1010_00110011101000___0011_001100111101100101;
		7'd58 : coef_acc =   57'b0011_11111111111111010___1010_00101011101100___0011_001111110110001100;
		7'd59 : coef_acc =   57'b0011_11111111111111010___1010_00100011110000___0011_010010101111110010;
		7'd60 : coef_acc =   57'b0011_11111111111111010___1010_00011011110100___0011_010101101010010111;
		7'd61 : coef_acc =   57'b0011_11111111111111010___1010_00010011111000___0011_011000100101111011;
		7'd62 : coef_acc =   57'b0011_11111111111111011___1010_00001011111100___0011_011011100010011110;
		7'd63 : coef_acc =   57'b0011_11111111111111011___1010_00000100000000___0011_011110100000000000;
		7'd64 : coef_acc =   57'b0011_11111111111111011___1001_11111100000100___0011_100001011110100001;
		7'd65 : coef_acc =   57'b0011_11111111111111011___1001_11110100001000___0011_100100011110000001;
		7'd66 : coef_acc =   57'b0011_11111111111111011___1001_11101100001100___0011_100111011110100000;
		7'd67 : coef_acc =   57'b0011_11111111111111011___1001_11100100010000___0011_101010011111111111;
		7'd68 : coef_acc =   57'b0011_11111111111111011___1001_11011100010100___0011_101101100010011100;
		7'd69 : coef_acc =   57'b0011_11111111111111011___1001_11010100011000___0011_110000100101111000;
		7'd70 : coef_acc =   57'b0011_11111111111111100___1001_11001100011100___0011_110011101010010011;
		7'd71 : coef_acc =   57'b0011_11111111111111100___1001_11000100011111___0011_110110101111101101;
		7'd72 : coef_acc =   57'b0011_11111111111111100___1001_10111100100011___0011_111001110110000110;
		7'd73 : coef_acc =   57'b0011_11111111111111100___1001_10110100100111___0011_111100111101011110;
		7'd74 : coef_acc =   57'b0011_11111111111111100___1001_10101100101011___0100_000000000101110101;
		7'd75 : coef_acc =   57'b0011_11111111111111100___1001_10100100101111___0100_000011001111001011;
		7'd76 : coef_acc =   57'b0011_11111111111111100___1001_10011100110011___0100_000110011001100001;
		7'd77 : coef_acc =   57'b0011_11111111111111100___1001_10010100110111___0100_001001100100110101;
		7'd78 : coef_acc =   57'b0011_11111111111111100___1001_10001100111011___0100_001100110001001000;
		7'd79 : coef_acc =   57'b0011_11111111111111100___1001_10000100111111___0100_001111111110011010;
		7'd80 : coef_acc =   57'b0011_11111111111111100___1001_01111101000011___0100_010011001100101011;
		7'd81 : coef_acc =   57'b0011_11111111111111100___1001_01110101000111___0100_010110011011111011;
		7'd82 : coef_acc =   57'b0011_11111111111111101___1001_01101101001011___0100_011001101100001010;
		7'd83 : coef_acc =   57'b0011_11111111111111101___1001_01100101001111___0100_011100111101011001;
		7'd84 : coef_acc =   57'b0011_11111111111111101___1001_01011101010011___0100_100000001111100110;
		7'd85 : coef_acc =   57'b0011_11111111111111101___1001_01010101010111___0100_100011100010110010;
		7'd86 : coef_acc =   57'b0011_11111111111111101___1001_01001101011011___0100_100110110110111101;
		7'd87 : coef_acc =   57'b0011_11111111111111101___1001_01000101011111___0100_101010001100000111;
		7'd88 : coef_acc =   57'b0011_11111111111111101___1001_00111101100011___0100_101101100010010001;
		7'd89 : coef_acc =   57'b0011_11111111111111101___1001_00110101100110___0100_110000111001011001;
		7'd90 : coef_acc =   57'b0011_11111111111111101___1001_00101101101010___0100_110100010001100000;
		7'd91 : coef_acc =   57'b0011_11111111111111101___1001_00100101101110___0100_110111101010100110;
		7'd92 : coef_acc =   57'b0011_11111111111111101___1001_00011101110010___0100_111011000100101011;
		7'd93 : coef_acc =   57'b0011_11111111111111101___1001_00010101110110___0100_111110011111110000;
		7'd94 : coef_acc =   57'b0011_11111111111111101___1001_00001101111010___0101_000001111011110011;
		7'd95 : coef_acc =   57'b0011_11111111111111101___1001_00000101111110___0101_000101011000110101;
		7'd96 : coef_acc =   57'b0011_11111111111111101___1000_11111110000010___0101_001000110110110110;
		7'd97 : coef_acc =   57'b0011_11111111111111101___1000_11110110000110___0101_001100010101110111;
		7'd98 : coef_acc =   57'b0011_11111111111111101___1000_11101110001010___0101_001111110101110110;
		7'd99 : coef_acc =   57'b0011_11111111111111101___1000_11100110001110___0101_010011010110110100;
		7'd100 : coef_acc =   57'b0011_11111111111111110___1000_11011110010010___0101_010110111000110010;
		7'd101 : coef_acc =   57'b0011_11111111111111110___1000_11010110010110___0101_011010011011101110;
		7'd102 : coef_acc =   57'b0011_11111111111111110___1000_11001110011010___0101_011101111111101001;
		7'd103 : coef_acc =   57'b0011_11111111111111110___1000_11000110011110___0101_100001100100100100;
		7'd104 : coef_acc =   57'b0011_11111111111111110___1000_10111110100010___0101_100101001010011101;
		7'd105 : coef_acc =   57'b0011_11111111111111110___1000_10110110100110___0101_101000110001010101;
		7'd106 : coef_acc =   57'b0011_11111111111111110___1000_10101110101010___0101_101100011001001101;
		7'd107 : coef_acc =   57'b0011_11111111111111110___1000_10100110101110___0101_110000000010000011;
		7'd108 : coef_acc =   57'b0011_11111111111111110___1000_10011110110010___0101_110011101011111000;
		7'd109 : coef_acc =   57'b0011_11111111111111110___1000_10010110110110___0101_110111010110101101;
		7'd110 : coef_acc =   57'b0011_11111111111111110___1000_10001110111010___0101_111011000010100000;
		7'd111 : coef_acc =   57'b0011_11111111111111110___1000_10000110111101___0101_111110101111010011;
		7'd112 : coef_acc =   57'b0011_11111111111111110___1000_01111111000001___0110_000010011101000100;
		7'd113 : coef_acc =   57'b0011_11111111111111110___1000_01110111000101___0110_000110001011110100;
		7'd114 : coef_acc =   57'b0011_11111111111111110___1000_01101111001001___0110_001001111011100100;
		7'd115 : coef_acc =   57'b0011_11111111111111110___1000_01100111001101___0110_001101101100010010;
		7'd116 : coef_acc =   57'b0011_11111111111111110___1000_01011111010001___0110_010001011110000000;
		7'd117 : coef_acc =   57'b0011_11111111111111110___1000_01010111010101___0110_010101010000101100;
		7'd118 : coef_acc =   57'b0011_11111111111111110___1000_01001111011001___0110_011001000100011000;
		7'd119 : coef_acc =   57'b0011_11111111111111110___1000_01000111011101___0110_011100111001000010;
		7'd120 : coef_acc =   57'b0011_11111111111111110___1000_00111111100001___0110_100000101110101100;
		7'd121 : coef_acc =   57'b0011_11111111111111110___1000_00110111100101___0110_100100100101010100;
		7'd122 : coef_acc =   57'b0011_11111111111111110___1000_00101111101001___0110_101000011100111100;
		7'd123 : coef_acc =   57'b0011_11111111111111110___1000_00100111101101___0110_101100010101100010;
		7'd124 : coef_acc =   57'b0011_11111111111111110___1000_00011111110001___0110_110000001111001000;
		7'd125 : coef_acc =   57'b0011_11111111111111110___1000_00010111110101___0110_110100001001101100;
		7'd126 : coef_acc =   57'b0011_11111111111111110___1000_00001111111001___0110_111000000101010000;
		7'd127 : coef_acc =   57'b0011_11111111111111110___1000_00000111111101___0110_111100000001110010;

endcase

always@(posedge clk)
	if(rst | ~en_coef)
		begin
			coef0<=21'd0;
			coef1<=18'd0;
			coef2<=18'd0;
		end
	else
		begin
			coef0<=coef_acc[20:0];
			coef1<=coef_acc[38:21];
		   coef2<=coef_acc[56:39];
		end

endmodule
