module ROM_coef(clk,rst,		// I: Global IO (clock, reset) 
			  en_coef,      // I: Module Enable signal
			  segment,    	// I: [6:0] Segment (Offset + ROM_trans)
			  coef0,        // O: [20:0] Coefficient 0
			  coef1,        // O: [17:0] Coefficient 1
			  coef2			// O: [17:0] Coefficient 2
			  );

input clk,rst;				// I: Global IO (clock, reset) 
input en_coef;      		// I: Module Enable signal
input [6:0]segment;    		// I: [6:0] Segment (Offset + ROM_trans)
output reg signed [20:0] coef0;	// O: [20:0] Coefficient 0
output reg signed [17:0] coef1;	// O: [17:0] Coefficient 1
output reg signed [17:0] coef2;	// O: [17:0] Coefficient 2

reg [56:0] coef_acc;

always@(*)
	case(segment)
		7'd   0 : coef_acc =   57'b1_11111110101100101___1011_11111010101100___001_000001101001110110;
		7'd   1 : coef_acc =   57'b1_11111111010110110___1011_11110001011100___001_000011110100111000;
		7'd   2 : coef_acc =   57'b1_11111111100100111___1011_11101001000011___001_000101111001110111;
		7'd   3 : coef_acc =   57'b1_11111111101011111___1011_11100000111001___001_000111111110000101;
		7'd   4 : coef_acc =   57'b1_11111111110000001___1011_11011000110101___001_001010000010100100;
		7'd   5 : coef_acc =   57'b1_11111111110010111___1011_11010000110011___001_001100000111101101;
		7'd   6 : coef_acc =   57'b1_11111111110100111___1011_11001000110011___001_001110001101100111;
		7'd   7 : coef_acc =   57'b1_11111111110110011___1011_11000000110100___001_010000010100011000;
		7'd   8 : coef_acc =   57'b1_11111111110111101___1011_10111000110110___001_010010011100000011;
		7'd   9 : coef_acc =   57'b1_11111111111000100___1011_10110000111000___001_010100100100101001;
		7'd  10 : coef_acc =   57'b1_11111111111001010___1011_10101000111010___001_010110101110001100;
		7'd  11 : coef_acc =   57'b1_11111111111001111___1011_10100000111101___001_011000111000101011;
		7'd  12 : coef_acc =   57'b1_11111111111010100___1011_10011001000000___001_011011000100001000;
		7'd  13 : coef_acc =   57'b1_11111111111010111___1011_10010001000011___001_011101010000100011;
		7'd  14 : coef_acc =   57'b1_11111111111011010___1011_10001001000110___001_011111011101111011;
		7'd  15 : coef_acc =   57'b1_11111111111011101___1011_10000001001001___001_100001101100010010;
		7'd  16 : coef_acc =   57'b1_11111111111100000___1011_01111001001101___001_100011111011100111;
		7'd  17 : coef_acc =   57'b1_11111111111100010___1011_01110001010000___001_100110001011111011;
		7'd  18 : coef_acc =   57'b1_11111111111100100___1011_01101001010100___001_101000011101001101;
		7'd  19 : coef_acc =   57'b1_11111111111100101___1011_01100001010111___001_101010101111011110;
		7'd  20 : coef_acc =   57'b1_11111111111100111___1011_01011001011011___001_101101000010101101;
		7'd  21 : coef_acc =   57'b1_11111111111101000___1011_01010001011110___001_101111010110111100;
		7'd  22 : coef_acc =   57'b1_11111111111101010___1011_01001001100010___001_110001101100001000;
		7'd  23 : coef_acc =   57'b1_11111111111101011___1011_01000001100110___001_110100000010010100;
		7'd  24 : coef_acc =   57'b1_11111111111101100___1011_00111001101001___001_110110011001011111;
		7'd  25 : coef_acc =   57'b1_11111111111101101___1011_00110001101101___001_111000110001101000;
		7'd  26 : coef_acc =   57'b1_11111111111101110___1011_00101001110001___001_111011001010110000;
		7'd  27 : coef_acc =   57'b1_11111111111101111___1011_00100001110100___001_111101100100111000;
		7'd  28 : coef_acc =   57'b1_11111111111101111___1011_00011001111000___001_111111111111111110;
		7'd  29 : coef_acc =   57'b1_11111111111110000___1011_00010001111100___010_000010011100000010;
		7'd  30 : coef_acc =   57'b1_11111111111110001___1011_00001010000000___010_000100111001000110;
		7'd  31 : coef_acc =   57'b1_11111111111110001___1011_00000010000100___010_000111010111001001;
		7'd  32 : coef_acc =   57'b1_11111111111110010___1010_11111010000111___010_001001110110001011;
		7'd  33 : coef_acc =   57'b1_11111111111110011___1010_11110010001011___010_001100010110001011;
		7'd  34 : coef_acc =   57'b1_11111111111110011___1010_11101010001111___010_001110110111001011;
		7'd  35 : coef_acc =   57'b1_11111111111110100___1010_11100010010011___010_010001011001001001;
		7'd  36 : coef_acc =   57'b1_11111111111110100___1010_11011010010111___010_010011111100000111;
		7'd  37 : coef_acc =   57'b1_11111111111110101___1010_11010010011011___010_010110100000000011;
		7'd  38 : coef_acc =   57'b1_11111111111110101___1010_11001010011110___010_011001000100111111;
		7'd  39 : coef_acc =   57'b1_11111111111110101___1010_11000010100010___010_011011101010111001;
		7'd  40 : coef_acc =   57'b1_11111111111110110___1010_10111010100110___010_011110010001110010;
		7'd  41 : coef_acc =   57'b1_11111111111110110___1010_10110010101010___010_100000111001101010;
		7'd  42 : coef_acc =   57'b1_11111111111110110___1010_10101010101110___010_100011100010100010;
		7'd  43 : coef_acc =   57'b1_11111111111110111___1010_10100010110010___010_100110001100011000;
		7'd  44 : coef_acc =   57'b1_11111111111110111___1010_10011010110110___010_101000110111001101;
		7'd  45 : coef_acc =   57'b1_11111111111110111___1010_10010010111010___010_101011100011000001;
		7'd  46 : coef_acc =   57'b1_11111111111111000___1010_10001010111101___010_101110001111110101;
		7'd  47 : coef_acc =   57'b1_11111111111111000___1010_10000011000001___010_110000111101100111;
		7'd  48 : coef_acc =   57'b1_11111111111111000___1010_01111011000101___010_110011101100011000;
		7'd  49 : coef_acc =   57'b1_11111111111111000___1010_01110011001001___010_110110011100001000;
		7'd  50 : coef_acc =   57'b1_11111111111111000___1010_01101011001101___010_111001001100110111;
		7'd  51 : coef_acc =   57'b1_11111111111111001___1010_01100011010001___010_111011111110100101;
		7'd  52 : coef_acc =   57'b1_11111111111111001___1010_01011011010101___010_111110110001010010;
		7'd  53 : coef_acc =   57'b1_11111111111111001___1010_01010011011001___011_000001100100111110;
		7'd  54 : coef_acc =   57'b1_11111111111111001___1010_01001011011101___011_000100011001101001;
		7'd  55 : coef_acc =   57'b1_11111111111111001___1010_01000011100001___011_000111001111010100;
		7'd  56 : coef_acc =   57'b1_11111111111111010___1010_00111011100101___011_001010000101111101;
		7'd  57 : coef_acc =   57'b1_11111111111111010___1010_00110011101000___011_001100111101100101;
		7'd  58 : coef_acc =   57'b1_11111111111111010___1010_00101011101100___011_001111110110001100;
		7'd  59 : coef_acc =   57'b1_11111111111111010___1010_00100011110000___011_010010101111110010;
		7'd  60 : coef_acc =   57'b1_11111111111111010___1010_00011011110100___011_010101101010010111;
		7'd  61 : coef_acc =   57'b1_11111111111111010___1010_00010011111000___011_011000100101111011;
		7'd  62 : coef_acc =   57'b1_11111111111111011___1010_00001011111100___011_011011100010011110;
		7'd  63 : coef_acc =   57'b1_11111111111111011___1010_00000100000000___011_011110100000000000;
		7'd  64 : coef_acc =   57'b1_11111111111111011___1001_11111100000100___011_100001011110100001;
		7'd  65 : coef_acc =   57'b1_11111111111111011___1001_11110100001000___011_100100011110000001;
		7'd  66 : coef_acc =   57'b1_11111111111111011___1001_11101100001100___011_100111011110100000;
		7'd  67 : coef_acc =   57'b1_11111111111111011___1001_11100100010000___011_101010011111111111;
		7'd  68 : coef_acc =   57'b1_11111111111111011___1001_11011100010100___011_101101100010011100;
		7'd  69 : coef_acc =   57'b1_11111111111111011___1001_11010100011000___011_110000100101111000;
		7'd  70 : coef_acc =   57'b1_11111111111111100___1001_11001100011100___011_110011101010010011;
		7'd  71 : coef_acc =   57'b1_11111111111111100___1001_11000100011111___011_110110101111101101;
		7'd  72 : coef_acc =   57'b1_11111111111111100___1001_10111100100011___011_111001110110000110;
		7'd  73 : coef_acc =   57'b1_11111111111111100___1001_10110100100111___011_111100111101011110;
		7'd  74 : coef_acc =   57'b1_11111111111111100___1001_10101100101011___100_000000000101110101;
		7'd  75 : coef_acc =   57'b1_11111111111111100___1001_10100100101111___100_000011001111001011;
		7'd  76 : coef_acc =   57'b1_11111111111111100___1001_10011100110011___100_000110011001100001;
		7'd  77 : coef_acc =   57'b1_11111111111111100___1001_10010100110111___100_001001100100110101;
		7'd  78 : coef_acc =   57'b1_11111111111111100___1001_10001100111011___100_001100110001001000;
		7'd  79 : coef_acc =   57'b1_11111111111111100___1001_10000100111111___100_001111111110011010;
		7'd  80 : coef_acc =   57'b1_11111111111111100___1001_01111101000011___100_010011001100101011;
		7'd  81 : coef_acc =   57'b1_11111111111111100___1001_01110101000111___100_010110011011111011;
		7'd  82 : coef_acc =   57'b1_11111111111111101___1001_01101101001011___100_011001101100001010;
		7'd  83 : coef_acc =   57'b1_11111111111111101___1001_01100101001111___100_011100111101011001;
		7'd  84 : coef_acc =   57'b1_11111111111111101___1001_01011101010011___100_100000001111100110;
		7'd  85 : coef_acc =   57'b1_11111111111111101___1001_01010101010111___100_100011100010110010;
		7'd  86 : coef_acc =   57'b1_11111111111111101___1001_01001101011011___100_100110110110111101;
		7'd  87 : coef_acc =   57'b1_11111111111111101___1001_01000101011111___100_101010001100000111;
		7'd  88 : coef_acc =   57'b1_11111111111111101___1001_00111101100011___100_101101100010010001;
		7'd  89 : coef_acc =   57'b1_11111111111111101___1001_00110101100110___100_110000111001011001;
		7'd  90 : coef_acc =   57'b1_11111111111111101___1001_00101101101010___100_110100010001100000;
		7'd  91 : coef_acc =   57'b1_11111111111111101___1001_00100101101110___100_110111101010100110;
		7'd  92 : coef_acc =   57'b1_11111111111111101___1001_00011101110010___100_111011000100101011;
		7'd  93 : coef_acc =   57'b1_11111111111111101___1001_00010101110110___100_111110011111110000;
		7'd  94 : coef_acc =   57'b1_11111111111111101___1001_00001101111010___101_000001111011110011;
		7'd  95 : coef_acc =   57'b1_11111111111111101___1001_00000101111110___101_000101011000110101;
		7'd  96 : coef_acc =   57'b1_11111111111111101___1000_11111110000010___101_001000110110110110;
		7'd  97 : coef_acc =   57'b1_11111111111111101___1000_11110110000110___101_001100010101110111;
		7'd  98 : coef_acc =   57'b1_11111111111111101___1000_11101110001010___101_001111110101110110;
		7'd  99 : coef_acc =   57'b1_11111111111111101___1000_11100110001110___101_010011010110110100;
		7'd 100 : coef_acc =   57'b1_11111111111111110___1000_11011110010010___101_010110111000110010;
		7'd 101 : coef_acc =   57'b1_11111111111111110___1000_11010110010110___101_011010011011101110;
		7'd 102 : coef_acc =   57'b1_11111111111111110___1000_11001110011010___101_011101111111101001;
		7'd 103 : coef_acc =   57'b1_11111111111111110___1000_11000110011110___101_100001100100100100;
		7'd 104 : coef_acc =   57'b1_11111111111111110___1000_10111110100010___101_100101001010011101;
		7'd 105 : coef_acc =   57'b1_11111111111111110___1000_10110110100110___101_101000110001010101;
		7'd 106 : coef_acc =   57'b1_11111111111111110___1000_10101110101010___101_101100011001001101;
		7'd 107 : coef_acc =   57'b1_11111111111111110___1000_10100110101110___101_110000000010000011;
		7'd 108 : coef_acc =   57'b1_11111111111111110___1000_10011110110010___101_110011101011111000;
		7'd 109 : coef_acc =   57'b1_11111111111111110___1000_10010110110110___101_110111010110101101;
		7'd 110 : coef_acc =   57'b1_11111111111111110___1000_10001110111010___101_111011000010100000;
		7'd 111 : coef_acc =   57'b1_11111111111111110___1000_10000110111101___101_111110101111010011;
		7'd 112 : coef_acc =   57'b1_11111111111111110___1000_01111111000001___110_000010011101000100;
		7'd 113 : coef_acc =   57'b1_11111111111111110___1000_01110111000101___110_000110001011110100;
		7'd 114 : coef_acc =   57'b1_11111111111111110___1000_01101111001001___110_001001111011100100;
		7'd 115 : coef_acc =   57'b1_11111111111111110___1000_01100111001101___110_001101101100010010;
		7'd 116 : coef_acc =   57'b1_11111111111111110___1000_01011111010001___110_010001011110000000;
		7'd 117 : coef_acc =   57'b1_11111111111111110___1000_01010111010101___110_010101010000101100;
		7'd 118 : coef_acc =   57'b1_11111111111111110___1000_01001111011001___110_011001000100011000;
		7'd 119 : coef_acc =   57'b1_11111111111111110___1000_01000111011101___110_011100111001000010;
		7'd 120 : coef_acc =   57'b1_11111111111111110___1000_00111111100001___110_100000101110101100;
		7'd 121 : coef_acc =   57'b1_11111111111111110___1000_00110111100101___110_100100100101010100;
		7'd 122 : coef_acc =   57'b1_11111111111111110___1000_00101111101001___110_101000011100111100;
		7'd 123 : coef_acc =   57'b1_11111111111111110___1000_00100111101101___110_101100010101100010;
		7'd 124 : coef_acc =   57'b1_11111111111111110___1000_00011111110001___110_110000001111001000;
		7'd 125 : coef_acc =   57'b1_11111111111111110___1000_00010111110101___110_110100001001101100;
		7'd 126 : coef_acc =   57'b1_11111111111111110___1000_00001111111001___110_111000000101010000;
		7'd 127 : coef_acc =   57'b1_11111111111111110___1000_00000111111101___110_111100000001110010;

endcase

always@(posedge clk)
	if(rst | ~en_coef)
		begin
			coef0<=21'd0;
			coef1<=18'd0;
			coef2<=18'd0;
		end
	else
		begin
			coef0<=coef_acc[20:0];
			coef1<=coef_acc[38:21];
		   coef2<=coef_acc[56:39];
		end

endmodule
